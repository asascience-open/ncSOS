netcdf timeSeriesProfile-Multidimensional-MultipeStations-H.5.1 {
dimensions:
	station = 2 ;
	profile = 4 ;
	z = 30 ;
	name_strlen = 50 ;
variables:
	double lat(station) ;
		lat:units = "degrees_north" ;
		lat:long_name = "station latitude" ;
		lat:standard_name = "latitude" ;
	double lon(station) ;
		lon:units = "degrees_east" ;
		lon:long_name = "station longitude" ;
		lon:standard_name = "longitude" ;
	int station_info(station) ;
		station_info:long_name = "station info" ;
	char station_name(station, name_strlen) ;
		station_name:cf_role = "timeseries_id" ;
		station_name:long_name = "station name" ;
	double alt(station, profile, z) ;
		alt:standard_name = "altitude" ;
		alt:long_name = "height above mean sea level" ;
		alt:units = "m" ;
		alt:positive = "up" ;
		alt:axis = "Z" ;
	int time(station, profile) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
	double temperature(station, profile, z) ;
		temperature:long_name = "Water Temperature" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:coordinates = "time lat lon alt" ;

// global attributes:
		:featureType = "timeSeriesProfile" ;
		:Conventions = "CF-1.6" ;
}
